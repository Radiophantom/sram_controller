
package sram_timings_pkg;

  parameter int TRC   = 45;
  parameter int TAA   = 45;
  parameter int TOHA  = 10;
  parameter int TDOE  = 22;
  parameter int TLZOE = 5;
  parameter int THZOE = 18;

  parameter int TWC   = 45;
  parameter int TAW   = 35;
  parameter int THA   = 0;
  parameter int TSA   = 0;
  parameter int TPWE  = 35;
  parameter int TSD   = 25;
  parameter int THD   = 0;
  parameter int THZWE = 18;
  parameter int TLZWE = 10;

endpackage

